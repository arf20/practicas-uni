//: version "2.0-b10etc2"
//: property encoding = "utf-8"
//: property locale = "es"
//: property prefix = "_GG"
//: property title = "sumador.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg [3:0] w8;    //: /sn:0 {0}(#:235,358)(#:235,409){1}
reg [3:0] w9;    //: /sn:0 {0}(#:388,367)(#:388,403){1}
wire w6;    //: /sn:0 {0}(265,269)(265,302)(239,302)(239,352){1}
wire w7;    //: /sn:0 {0}(300,269)(300,331)(249,331)(249,352){1}
wire w14;    //: /sn:0 {0}(303,37)(303,70)(475,70)(475,107){1}
wire w15;    //: /sn:0 {0}(293,37)(293,86)(411,86)(411,107){1}
wire w4;    //: /sn:0 {0}(194,269)(194,337)(219,337)(219,352){1}
wire w0;    //: /sn:0 {0}(372,361)(372,342)(347,342)(347,269){1}
wire w3;    //: /sn:0 {0}(471,269)(471,346)(402,346)(402,361){1}
wire w1;    //: /sn:0 {0}(382,361)(382,284)(381,284)(381,269){1}
wire w18;    //: /sn:0 {0}(212,107)(212,47)(273,47)(273,37){1}
wire w17;    //: /sn:0 {0}(283,37)(283,95)(287,95)(287,107){1}
wire w2;    //: /sn:0 {0}(392,361)(392,284)(425,284)(425,269){1}
wire w12;    //: /sn:0 {0}(243,-24)(243,4)(155,4)(155,193)(176,193){1}
wire [3:0] w13;    //: /sn:0 {0}(#:288,31)(288,2)(289,2)(289,-15){1}
wire w5;    //: /sn:0 {0}(229,269)(229,352){1}
//: enddecls

  //: DIP g4 (w8) @(235,420) /sn:0 /R:2 /w:[ 1 ] /st:0 /dn:1
  //: LED g3 (w12) @(243,-31) /sn:0 /w:[ 0 ] /type:0
  assign w13 = {w18, w17, w15, w14}; //: CONCAT g2  @(288,32) /sn:0 /R:1 /w:[ 0 1 0 0 0 ] /dr:0 /tp:0 /drp:1
  //: LED g1 (w13) @(289,-22) /sn:0 /w:[ 1 ] /type:2
  //: DIP g6 (w9) @(388,414) /sn:0 /R:2 /w:[ 1 ] /st:0 /dn:1
  assign {w0, w1, w2, w3} = w9; //: CONCAT g7  @(387,366) /sn:0 /R:3 /w:[ 0 0 0 1 0 ] /dr:1 /tp:0 /drp:0
  assign {w4, w5, w6, w7} = w8; //: CONCAT g5  @(234,357) /sn:0 /R:3 /w:[ 1 1 1 1 0 ] /dr:1 /tp:0 /drp:0
  sumador4bits g0 (.a0(w7), .a1(w6), .a2(w5), .a3(w4), .b0(w3), .b1(w2), .b2(w1), .b3(w0), .r0(w14), .r1(w15), .r2(w17), .r3(w18), .cout(w12));   //: @(177, 108) /sz:(320, 160) /sn:0 /p:[ Bi0>0 Bi1>0 Bi2>0 Bi3>0 Bi4>0 Bi5>1 Bi6>1 Bi7>1 To0<1 To1<1 To2<1 To3<0 Lo0<1 ]

endmodule
//: /netlistEnd

//: /netlistBegin sumador4bits
module sumador4bits(r3, a3, a1, b2, a0, r1, r2, cout, b1, b3, r0, b0, a2);
//: interface  /sz:(320, 160) /bd:[ Bi0>a0(123/320) Bi1>a1(88/320) Bi2>a2(52/320) Bi3>a3(17/320) Bi4>b0(294/320) Bi5>b1(248/320) Bi6>b2(204/320) Bi7>b3(170/320) To0<r0(298/320) To1<r1(234/320) To2<r2(110/320) To3<r3(35/320) Lo0<cout(85/160) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input a2;    //: /sn:0 {0}(312,263)(312,316){1}
input b2;    //: /sn:0 {0}(352,263)(352,294)(354,294)(354,309){1}
input a3;    //: /sn:0 {0}(156,263)(156,293)(155,293)(155,308){1}
input b3;    //: /sn:0 {0}(196,263)(196,296)(195,296)(195,302){1}
output r1;    //: /sn:0 {0}(461,123)(461,150)(462,150)(462,165){1}
output r3;    //: /sn:0 {0}(155,121)(155,150)(156,150)(156,165){1}
input a1;    //: /sn:0 {0}(462,263)(462,314){1}
output r0;    //: /sn:0 {0}(611,117)(611,165){1}
input b1;    //: /sn:0 {0}(503,311)(503,286)(502,286)(502,263){1}
input a0;    //: /sn:0 {0}(611,263)(611,316){1}
input b0;    //: /sn:0 {0}(651,263)(651,309)(654,309)(654,318){1}
output cout;    //: /sn:0 {0}(70,184)(120,184)(120,182)(135,182){1}
supply0 w9;    //: /sn:0 {0}(680,182)(725,182)(725,211){1}
output r2;    //: /sn:0 {0}(312,122)(312,165){1}
wire w7;    //: /sn:0 {0}(381,182)(441,182){1}
wire w12;    //: /sn:0 {0}(531,182)(590,182){1}
wire w2;    //: /sn:0 {0}(225,182)(291,182){1}
//: enddecls

  //: GROUND g4 (w9) @(725,217) /sn:0 /w:[ 1 ]
  //: OUT g8 (r3) @(155,124) /sn:0 /R:1 /w:[ 0 ]
  sumador g3 (.a(a0), .b(b0), .c(w9), .r(r0), .ci(w12));   //: @(591, 166) /sz:(88, 96) /sn:0 /p:[ Bi0>0 Bi1>0 Ri0>0 To0<1 Lo0<1 ]
  //: IN g13 (a3) @(155,310) /sn:0 /R:1 /w:[ 1 ]
  sumador g2 (.a(a1), .b(b1), .c(w12), .r(r1), .ci(w7));   //: @(442, 166) /sz:(88, 96) /sn:0 /p:[ Bi0>0 Bi1>1 Ri0>0 To0<1 Lo0<1 ]
  sumador g1 (.a(a2), .b(b2), .c(w7), .r(r2), .ci(w2));   //: @(292, 166) /sz:(88, 96) /sn:0 /p:[ Bi0>0 Bi1>0 Ri0>0 To0<1 Lo0<1 ]
  //: IN g11 (a1) @(462,316) /sn:0 /R:1 /w:[ 1 ]
  //: IN g16 (b2) @(354,311) /sn:0 /R:1 /w:[ 1 ]
  //: IN g10 (a0) @(611,318) /sn:0 /R:1 /w:[ 1 ]
  //: OUT g6 (r1) @(461,126) /sn:0 /R:1 /w:[ 0 ]
  //: OUT g7 (r2) @(312,125) /sn:0 /R:1 /w:[ 0 ]
  //: OUT g9 (cout) @(73,184) /sn:0 /R:2 /w:[ 0 ]
  //: IN g15 (b1) @(503,313) /sn:0 /R:1 /w:[ 0 ]
  //: IN g17 (b3) @(195,304) /sn:0 /R:1 /w:[ 1 ]
  //: OUT g5 (r0) @(611,120) /sn:0 /R:1 /w:[ 0 ]
  //: IN g14 (b0) @(654,320) /sn:0 /R:1 /w:[ 1 ]
  sumador g0 (.a(a3), .b(b3), .c(w2), .r(r3), .ci(cout));   //: @(136, 166) /sz:(88, 96) /sn:0 /p:[ Bi0>0 Bi1>0 Ri0>0 To0<1 Lo0<1 ]
  //: IN g12 (a2) @(312,318) /sn:0 /R:1 /w:[ 1 ]

endmodule
//: /netlistEnd

//: /netlistBegin sumador
module sumador(a, c, ci, r, b);
//: interface  /sz:(40, 40) /bd:[ ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input b;    //: /sn:0 {0}(130,167)(130,190)(129,190)(129,228){1}
//: {2}(131,230)(265,230)(265,198){3}
//: {4}(129,232)(129,260){5}
output r;    //: /sn:0 {0}(125,53)(125,110)(129,110)(129,125){1}
output ci;    //: /sn:0 {0}(245,49)(245,93)(249,93)(249,108){1}
input a;    //: /sn:0 {0}(98,167)(98,212){1}
//: {2}(100,214)(249,214)(249,198){3}
//: {4}(98,216)(98,265){5}
input c;    //: /sn:0 {0}(157,261)(157,250){1}
//: {2}(159,248)(281,248)(281,198){3}
//: {4}(157,246)(157,180)(158,180)(158,167){5}
//: enddecls

  //: IN g4 (a) @(98,267) /sn:0 /R:1 /w:[ 5 ]
  //: IN g8 (c) @(157,263) /sn:0 /R:1 /w:[ 0 ]
  //: OUT g3 (ci) @(245,52) /sn:0 /R:1 /w:[ 0 ]
  //: OUT g2 (r) @(125,56) /sn:0 /R:1 /w:[ 0 ]
  acarreo g1 (.a(a), .b(b), .c(c), .ci(ci));   //: @(233, 109) /sz:(64, 88) /R:1 /sn:0 /p:[ Bi0>3 Bi1>3 Bi2>3 To0<1 ]
  //: IN g6 (b) @(129,262) /sn:0 /R:1 /w:[ 5 ]
  //: joint g7 (b) @(129, 230) /w:[ 2 1 -1 4 ]
  //: joint g9 (c) @(157, 248) /w:[ 2 4 -1 1 ]
  //: joint g5 (a) @(98, 214) /w:[ 2 1 -1 4 ]
  resultado g0 (.a(a), .b(b), .c(c), .r(r));   //: @(87, 126) /sz:(92, 40) /sn:0 /p:[ Bi0>0 Bi1>0 Bi2>5 To0<1 ]

endmodule
//: /netlistEnd

//: /netlistBegin resultado
module resultado(b, a, c, r);
//: interface  /sz:(40, 40) /bd:[ ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input b;    //: /sn:0 {0}(91,174)(91,228)(144,228){1}
//: {2}(148,228)(175,228){3}
//: {4}(179,228)(213,228)(213,174){5}
//: {6}(177,226)(177,216)(172,216)(172,174){7}
//: {8}(146,226)(146,216)(127,216)(127,174){9}
//: {10}(146,230)(146,256){11}
output r;    //: /sn:0 {0}(156,53)(156,71){1}
input a;    //: /sn:0 {0}(92,258)(92,244){1}
//: {2}(94,242)(104,242)(104,241)(120,241){3}
//: {4}(124,241)(142,241)(142,242)(165,242){5}
//: {6}(169,242)(208,242)(208,174){7}
//: {8}(167,240)(167,174){9}
//: {10}(122,239)(122,174){11}
//: {12}(90,242)(86,242)(86,174){13}
input c;    //: /sn:0 {0}(218,174)(218,187)(235,187)(235,201)(228,201){1}
//: {2}(224,201)(178,201){3}
//: {4}(176,199)(176,189)(177,189)(177,174){5}
//: {6}(174,201)(133,201){7}
//: {8}(131,199)(131,189)(132,189)(132,174){9}
//: {10}(129,201)(96,201)(96,174){11}
//: {12}(226,203)(226,258){13}
wire w0;    //: /sn:0 {0}(91,153)(91,139)(122,139)(122,108)(149,108)(149,92){1}
wire w1;    //: /sn:0 {0}(154,92)(154,125)(127,125)(127,153){1}
wire w18;    //: /sn:0 {0}(159,92)(159,112)(172,112)(172,153){1}
wire w13;    //: /sn:0 {0}(213,153)(213,92)(164,92)(164,92){1}
//: enddecls

  _GGAND3 #(8) g4 (.I0(a), .I1(!b), .I2(!c), .Z(w18));   //: @(172,163) /sn:0 /R:1 /w:[ 9 7 5 1 ]
  //: IN g8 (b) @(146,258) /sn:0 /R:1 /w:[ 11 ]
  _GGAND3 #(8) g3 (.I0(!a), .I1(b), .I2(!c), .Z(w1));   //: @(127,163) /sn:0 /R:1 /w:[ 11 9 9 1 ]
  //: joint g13 (b) @(177, 228) /w:[ 4 6 3 -1 ]
  _GGAND3 #(8) g2 (.I0(!a), .I1(!b), .I2(c), .Z(w0));   //: @(91,163) /sn:0 /R:1 /w:[ 13 0 11 0 ]
  _GGOR4 #(10) g1 (.I0(w0), .I1(w1), .I2(w18), .I3(w13), .Z(r));   //: @(156,81) /sn:0 /R:1 /w:[ 1 0 0 1 1 ]
  //: joint g11 (a) @(167, 242) /w:[ 6 8 5 -1 ]
  //: joint g16 (c) @(226, 201) /w:[ 1 -1 2 12 ]
  //: joint g10 (a) @(122, 241) /w:[ 4 10 3 -1 ]
  //: IN g6 (a) @(92,260) /sn:0 /R:1 /w:[ 0 ]
  //: IN g7 (c) @(226,260) /sn:0 /R:1 /w:[ 13 ]
  //: joint g9 (a) @(92, 242) /w:[ 2 -1 12 1 ]
  //: joint g15 (c) @(176, 201) /w:[ 3 4 6 -1 ]
  _GGAND3 #(8) g5 (.I0(a), .I1(b), .I2(c), .Z(w13));   //: @(213,163) /sn:0 /R:1 /w:[ 7 5 0 0 ]
  //: joint g14 (c) @(131, 201) /w:[ 7 8 10 -1 ]
  //: OUT g0 (r) @(156,56) /sn:0 /R:1 /w:[ 0 ]
  //: joint g12 (b) @(146, 228) /w:[ 2 8 1 10 ]

endmodule
//: /netlistEnd

//: /netlistBegin acarreo
module acarreo(b, c, a, ci);
//: interface  /sz:(40, 40) /bd:[ ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input b;    //: /sn:0 {0}(102,185)(102,228)(174,228){1}
//: {2}(178,228)(218,228)(218,183){3}
//: {4}(176,230)(176,259){5}
output ci;    //: /sn:0 {0}(161,29)(161,78){1}
input a;    //: /sn:0 {0}(89,259)(89,243){1}
//: {2}(91,241)(158,241)(158,185){3}
//: {4}(89,239)(89,198)(97,198)(97,185){5}
input c;    //: /sn:0 {0}(163,185)(163,209)(221,209){1}
//: {2}(223,207)(223,183){3}
//: {4}(223,211)(223,266){5}
wire w0;    //: /sn:0 {0}(156,99)(156,127)(100,127)(100,164){1}
wire w3;    //: /sn:0 {0}(166,99)(166,147)(221,147)(221,162){1}
wire w1;    //: /sn:0 {0}(161,99)(161,164){1}
//: enddecls

  _GGAND2 #(6) g4 (.I0(b), .I1(c), .Z(w3));   //: @(221,172) /sn:0 /R:1 /w:[ 3 3 1 ]
  //: joint g8 (a) @(89, 241) /w:[ 2 4 -1 1 ]
  _GGAND2 #(6) g3 (.I0(a), .I1(c), .Z(w1));   //: @(161,174) /sn:0 /R:1 /w:[ 3 0 1 ]
  _GGAND2 #(6) g2 (.I0(a), .I1(b), .Z(w0));   //: @(100,174) /sn:0 /R:1 /w:[ 5 0 1 ]
  _GGOR3 #(8) g1 (.I0(w0), .I1(w1), .I2(w3), .Z(ci));   //: @(161,88) /sn:0 /R:1 /w:[ 0 0 0 1 ]
  //: joint g10 (c) @(223, 209) /w:[ -1 2 1 4 ]
  //: IN g6 (b) @(176,261) /sn:0 /R:1 /w:[ 5 ]
  //: IN g7 (c) @(223,268) /sn:0 /R:1 /w:[ 5 ]
  //: joint g9 (b) @(176, 228) /w:[ 2 -1 1 4 ]
  //: IN g5 (a) @(89,261) /sn:0 /R:1 /w:[ 0 ]
  //: OUT g0 (ci) @(161,32) /sn:0 /R:1 /w:[ 0 ]

endmodule
//: /netlistEnd

