//: version "2.0-b10etc2"
//: property encoding = "utf-8"
//: property locale = "es"
//: property prefix = "_GG"
//: property title = "PANIC.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg [3:0] w5;    //: /sn:0 {0}(#:542,43)(#:542,101){1}
wire w32;    //: /sn:0 {0}(12,481)(99,481)(99,482)(236,482){1}
//: {2}(240,482)(253,482){3}
//: {4}(238,480)(238,464){5}
//: {6}(240,462)(253,462){7}
//: {8}(238,460)(238,444){9}
//: {10}(240,442)(253,442){11}
//: {12}(238,440)(238,422)(253,422){13}
wire w6;    //: /sn:0 {0}(164,264)(164,567){1}
//: {2}(166,569)(746,569){3}
//: {4}(748,567)(748,531){5}
//: {6}(748,527)(748,410){7}
//: {8}(748,406)(748,186){9}
//: {10}(748,182)(748,72)(638,72)(638,33){11}
//: {12}(746,184)(552,184){13}
//: {14}(550,182)(550,112){15}
//: {16}(548,184)(456,184)(456,185)(368,185){17}
//: {18}(550,186)(550,196)(546,196)(546,199){19}
//: {20}(746,408)(736,408)(736,409)(592,409){21}
//: {22}(746,529)(539,529){23}
//: {24}(748,571)(748,700)(399,700){25}
//: {26}(162,569)(-9,569)(-9,546){27}
wire w14;    //: /sn:0 {0}(360,331)(375,331)(375,349){1}
//: {2}(377,351)(391,351)(391,246)(405,246){3}
//: {4}(373,351)(360,351){5}
//: {6}(375,353)(375,369){7}
//: {8}(373,371)(360,371){9}
//: {10}(375,373)(375,391)(360,391){11}
wire w16;    //: /sn:0 {0}(316,635)(316,520){1}
//: {2}(318,518)(336,518)(336,503){3}
//: {4}(316,516)(316,503){5}
//: {6}(314,518)(298,518){7}
//: {8}(296,516)(296,503){9}
//: {10}(294,518)(276,518)(276,503){11}
wire w4;    //: /sn:0 {0}(276,305)(276,290)(294,290){1}
//: {2}(298,290)(314,290){3}
//: {4}(318,290)(336,290)(336,305){5}
//: {6}(316,288)(316,210)(315,210)(315,202){7}
//: {8}(316,292)(316,305){9}
//: {10}(296,292)(296,305){11}
wire w3;    //: /sn:0 {0}(44,264)(44,622){1}
//: {2}(46,624)(443,624)(443,625)(641,625){3}
//: {4}(643,623)(643,483){5}
//: {6}(643,479)(643,362){7}
//: {8}(643,358)(643,138){9}
//: {10}(645,136)(655,136)(655,56)(752,56)(752,32){11}
//: {12}(641,136)(522,136){13}
//: {14}(520,134)(520,112){15}
//: {16}(518,136)(428,136){17}
//: {18}(424,136)(394,136)(394,137)(368,137){19}
//: {20}(426,138)(426,199){21}
//: {22}(641,360)(631,360)(631,361)(592,361){23}
//: {24}(641,481)(539,481){25}
//: {26}(643,627)(643,652)(399,652){27}
//: {28}(42,624)(-129,624)(-129,546){29}
wire w0;    //: /sn:0 {0}(124,264)(124,583){1}
//: {2}(126,585)(714,585){3}
//: {4}(716,583)(716,515){5}
//: {6}(716,511)(716,395){7}
//: {8}(716,391)(716,170){9}
//: {10}(716,166)(716,121)(703,121)(703,84)(678,84)(678,32){11}
//: {12}(714,168)(542,168){13}
//: {14}(540,166)(540,112){15}
//: {16}(538,168)(508,168){17}
//: {18}(504,168)(434,168)(434,169)(368,169){19}
//: {20}(506,170)(506,199){21}
//: {22}(714,393)(592,393){23}
//: {24}(714,513)(539,513){25}
//: {26}(716,587)(716,684)(399,684){27}
//: {28}(122,585)(-49,585)(-49,546){29}
wire w21;    //: /sn:0 {0}(360,420)(375,420)(375,438){1}
//: {2}(373,440)(360,440){3}
//: {4}(375,442)(375,458){5}
//: {6}(373,460)(360,460){7}
//: {8}(375,462)(375,478){9}
//: {10}(373,480)(360,480){11}
//: {12}(375,482)(375,492)(374,492)(374,481)(435,481){13}
wire w28;    //: /sn:0 {0}(185,242)(210,242)(210,326)(234,326){1}
//: {2}(238,326)(253,326){3}
//: {4}(236,328)(236,344){5}
//: {6}(238,346)(253,346){7}
//: {8}(236,348)(236,364){9}
//: {10}(238,366)(253,366){11}
//: {12}(236,368)(236,386)(253,386){13}
wire w12;    //: /sn:0 {0}(276,397)(276,382)(294,382){1}
//: {2}(298,382)(314,382){3}
//: {4}(318,382)(334,382){5}
//: {6}(336,380)(336,361)(488,361){7}
//: {8}(336,384)(336,397){9}
//: {10}(316,384)(316,397){11}
//: {12}(296,384)(296,397){13}
wire w2;    //: /sn:0 {0}(84,264)(84,602){1}
//: {2}(86,604)(678,604){3}
//: {4}(680,602)(680,499){5}
//: {6}(680,495)(680,378){7}
//: {8}(680,374)(680,154){9}
//: {10}(680,150)(680,108)(716,108)(716,32){11}
//: {12}(678,152)(532,152){13}
//: {14}(530,150)(530,112){15}
//: {16}(528,152)(469,152){17}
//: {18}(465,152)(415,152)(415,153)(368,153){19}
//: {20}(467,154)(467,178)(466,178)(466,199){21}
//: {22}(678,376)(668,376)(668,377)(592,377){23}
//: {24}(678,497)(539,497){25}
//: {26}(680,606)(680,668)(399,668){27}
//: {28}(82,604)(-89,604)(-89,546){29}
//: enddecls

  segmentoF g61 (.a0(w3), .a1(w2), .a2(w0), .a3(w6), .E(w28));   //: @(24, 183) /sz:(160, 80) /sn:0 /p:[ Bi0>0 Bi1>0 Bi2>0 Bi3>0 Ro0<0 ]
  //: LED g8 (w12) @(276,404) /sn:0 /R:2 /w:[ 0 ] /type:0
  //: LED g4 (w4) @(336,312) /sn:0 /R:2 /w:[ 5 ] /type:0
  //: joint g58 (w0) @(716, 585) /w:[ -1 4 3 26 ]
  //: joint g55 (w0) @(716, 513) /w:[ -1 6 24 5 ]
  //: joint g37 (w2) @(467, 152) /w:[ 17 -1 18 20 ]
  //: LED g13 (w14) @(353,391) /sn:0 /R:1 /w:[ 11 ] /type:0
  //: LED g3 (w4) @(316,312) /sn:0 /R:2 /w:[ 9 ] /type:0
  //: joint g34 (w14) @(375, 351) /w:[ 2 1 4 6 ]
  //: joint g51 (w32) @(238, 442) /w:[ 10 12 -1 9 ]
  //: LED g76 (w3) @(752,25) /sn:0 /w:[ 11 ] /type:0
  //: joint g65 (w21) @(375, 480) /w:[ -1 9 10 12 ]
  //: LED g2 (w4) @(296,312) /sn:0 /R:2 /w:[ 11 ] /type:0
  //: joint g77 (w12) @(336, 382) /w:[ -1 6 5 8 ]
  //: joint g59 (w12) @(296, 382) /w:[ 2 -1 1 12 ]
  //: LED g1 (w4) @(276,312) /sn:0 /R:2 /w:[ 0 ] /type:0
  segmentoG g72 (.a0(w3), .a1(w2), .a2(w0), .a3(w6), .G(w12));   //: @(489, 345) /sz:(102, 96) /sn:0 /p:[ Ri0>23 Ri1>23 Ri2>23 Ri3>21 Lo0<7 ]
  //: joint g64 (w28) @(236, 366) /w:[ 10 9 -1 12 ]
  //: LED g16 (w14) @(353,331) /sn:0 /R:1 /w:[ 0 ] /type:0
  //: LED g11 (w16) @(316,496) /sn:0 /w:[ 5 ] /type:0
  //: joint g50 (w2) @(680, 497) /w:[ -1 6 24 5 ]
  //: LED g28 (w32) @(260,482) /sn:0 /R:3 /w:[ 3 ] /type:0
  //: LED g10 (w16) @(296,496) /sn:0 /w:[ 9 ] /type:0
  //: joint g78 (w3) @(643, 360) /w:[ -1 8 22 7 ]
  assign {w6, w0, w2, w3} = w5; //: CONCAT g32  @(535,107) /sn:0 /R:1 /w:[ 15 15 15 15 1 ] /dr:1 /tp:0 /drp:0
  //: LED g27 (w32) @(260,462) /sn:0 /R:3 /w:[ 7 ] /type:0
  //: LED g19 (w21) @(353,440) /sn:0 /R:1 /w:[ 3 ] /type:0
  //: joint g69 (w0) @(124, 585) /w:[ 2 1 28 -1 ]
  //: joint g38 (w3) @(426, 136) /w:[ 17 -1 18 20 ]
  //: LED g6 (w12) @(316,404) /sn:0 /R:2 /w:[ 11 ] /type:0
  //: LED g75 (w2) @(716,25) /sn:0 /w:[ 11 ] /type:0
  //: joint g57 (w6) @(748, 569) /w:[ -1 4 3 24 ]
  //: LED g9 (w16) @(276,496) /sn:0 /w:[ 11 ] /type:0
  //: LED g7 (w12) @(296,404) /sn:0 /R:2 /w:[ 13 ] /type:0
  segmentoE g53 (.a0(w3), .a1(w2), .a2(w0), .a3(w6), .E(w32));   //: @(-149, 465) /sz:(160, 80) /sn:0 /p:[ Bi0>29 Bi1>29 Bi2>29 Bi3>27 Ro0<0 ]
  //: joint g71 (w3) @(44, 624) /w:[ 2 1 28 -1 ]
  //: DIP g31 (w5) @(542,33) /sn:0 /w:[ 0 ] /st:15 /dn:1
  //: LED g20 (w21) @(353,460) /sn:0 /R:1 /w:[ 7 ] /type:0
  //: LED g15 (w14) @(353,351) /sn:0 /R:1 /w:[ 5 ] /type:0
  //: joint g68 (w6) @(164, 569) /w:[ 2 1 26 -1 ]
  //: joint g67 (w3) @(643, 625) /w:[ -1 4 3 26 ]
  segmentoC g39 (.a0(w3), .a1(w2), .a2(w0), .a3(w6), .C(w21));   //: @(436, 465) /sz:(102, 96) /sn:0 /p:[ Ri0>25 Ri1>25 Ri2>25 Ri3>23 Lo0<13 ]
  //: joint g48 (w0) @(540, 168) /w:[ 13 14 16 -1 ]
  //: joint g43 (w3) @(520, 136) /w:[ 13 14 16 -1 ]
  //: LED g73 (w6) @(638,26) /sn:0 /w:[ 11 ] /type:0
  //: joint g62 (w28) @(236, 326) /w:[ 2 -1 1 4 ]
  //: joint g29 (w4) @(296, 290) /w:[ 2 -1 1 10 ]
  //: LED g25 (w32) @(260,422) /sn:0 /R:3 /w:[ 13 ] /type:0
  //: LED g17 (w21) @(353,480) /sn:0 /R:1 /w:[ 11 ] /type:0
  //: joint g63 (w28) @(236, 346) /w:[ 6 5 -1 8 ]
  //: joint g42 (w21) @(375, 460) /w:[ -1 5 6 8 ]
  //: joint g52 (w32) @(238, 462) /w:[ 6 8 -1 5 ]
  //: joint g83 (w0) @(716, 168) /w:[ -1 10 12 9 ]
  //: LED g74 (w0) @(678,25) /sn:0 /w:[ 11 ] /type:0
  //: joint g56 (w6) @(748, 529) /w:[ -1 6 22 5 ]
  //: LED g14 (w14) @(353,371) /sn:0 /R:1 /w:[ 9 ] /type:0
  //: LED g5 (w12) @(336,404) /sn:0 /R:2 /w:[ 9 ] /type:0
  //: joint g47 (w2) @(530, 152) /w:[ 13 14 16 -1 ]
  //: joint g44 (w16) @(296, 518) /w:[ 7 8 10 -1 ]
  //: joint g79 (w2) @(680, 376) /w:[ -1 8 22 7 ]
  //: joint g80 (w0) @(716, 393) /w:[ -1 8 22 7 ]
  //: joint g85 (w3) @(643, 136) /w:[ 10 -1 12 9 ]
  //: joint g84 (w2) @(680, 152) /w:[ -1 10 12 9 ]
  //: joint g36 (w0) @(506, 168) /w:[ 17 -1 18 20 ]
  //: LED g24 (w28) @(260,346) /sn:0 /R:3 /w:[ 7 ] /type:0
  //: LED g21 (w28) @(260,326) /sn:0 /R:3 /w:[ 3 ] /type:0
  //: LED g23 (w28) @(260,366) /sn:0 /R:3 /w:[ 11 ] /type:0
  //: joint g41 (w21) @(375, 440) /w:[ -1 1 2 4 ]
  //: joint g81 (w6) @(748, 184) /w:[ -1 10 12 9 ]
  segmentoB g40 (.a0(w3), .a1(w2), .a2(w0), .a3(w6), .B(w14));   //: @(406, 200) /sz:(160, 96) /sn:0 /p:[ Ti0>21 Ti1>21 Ti2>21 Ti3>19 Lo0<3 ]
  //: joint g54 (w32) @(238, 482) /w:[ 2 4 1 -1 ]
  //: joint g60 (w12) @(316, 382) /w:[ 4 -1 3 10 ]
  //: joint g70 (w2) @(84, 604) /w:[ 2 1 28 -1 ]
  //: LED g26 (w32) @(260,442) /sn:0 /R:3 /w:[ 11 ] /type:0
  //: LED g22 (w28) @(260,386) /sn:0 /R:3 /w:[ 13 ] /type:0
  segmentoA g0 (.A0(w3), .A1(w2), .A2(w0), .A3(w6), .A(w4));   //: @(265, 121) /sz:(102, 80) /sn:0 /p:[ Ri0>19 Ri1>19 Ri2>19 Ri3>17 Bo0<7 ]
  //: joint g35 (w14) @(375, 371) /w:[ -1 7 8 10 ]
  //: joint g45 (w16) @(316, 518) /w:[ 2 4 6 1 ]
  segmentoD g46 (.a0(w3), .a1(w2), .a2(w0), .a3(w6), .D(w16));   //: @(296, 636) /sz:(102, 80) /sn:0 /p:[ Ri0>27 Ri1>27 Ri2>27 Ri3>25 To0<0 ]
  //: joint g66 (w2) @(680, 604) /w:[ -1 4 3 26 ]
  //: joint g82 (w6) @(748, 408) /w:[ -1 8 20 7 ]
  //: LED g18 (w21) @(353,420) /sn:0 /R:1 /w:[ 0 ] /type:0
  //: LED g12 (w16) @(336,496) /sn:0 /w:[ 3 ] /type:0
  //: joint g33 (w6) @(550, 184) /w:[ 13 14 16 18 ]
  //: joint g30 (w4) @(316, 290) /w:[ 4 6 3 8 ]
  //: joint g49 (w3) @(643, 481) /w:[ -1 6 24 5 ]

endmodule
//: /netlistEnd

//: /netlistBegin segmentoA
module segmentoA(A2, A0, A3, A1, A);
//: interface  /sz:(102, 80) /bd:[ Ri0>A3(64/80) Ri1>A2(48/80) Ri2>A1(32/80) Ri3>A0(16/80) Bo0<A(50/102) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input A0;    //: /sn:0 {0}(351,281)(351,319)(36,319){1}
//: {2}(32,319)(5,319){3}
//: {4}(34,321)(34,337)(49,337){5}
input A3;    //: /sn:0 {0}(216,286)(216,415)(34,415){1}
//: {2}(30,415)(5,415){3}
//: {4}(32,417)(32,444)(49,444){5}
output A;    //: /sn:0 {0}(214,88)(214,156)(219,156)(219,171){1}
input A2;    //: /sn:0 {0}(5,386)(32,386){1}
//: {2}(36,386)(346,386)(346,281){3}
//: {4}(34,388)(34,399)(49,399){5}
input A1;    //: /sn:0 {0}(149,286)(149,353){1}
//: {2}(151,355)(286,355)(286,284){3}
//: {4}(147,355)(5,355){5}
wire w7;    //: /sn:0 {0}(65,399)(79,399){1}
//: {2}(83,399)(221,399)(221,286){3}
//: {4}(81,397)(81,287){5}
wire w14;    //: /sn:0 {0}(229,192)(229,204)(346,204)(346,260){1}
wire w1;    //: /sn:0 {0}(65,337)(84,337){1}
//: {2}(88,337)(154,337)(154,286){3}
//: {4}(86,335)(86,287){5}
wire w8;    //: /sn:0 {0}(219,265)(219,192){1}
wire w11;    //: /sn:0 {0}(224,192)(224,248)(284,248)(284,263){1}
wire w2;    //: /sn:0 {0}(209,192)(209,209)(84,209)(84,266){1}
wire w5;    //: /sn:0 {0}(214,192)(214,250)(152,250)(152,265){1}
wire w9;    //: /sn:0 {0}(281,284)(281,442){1}
//: {2}(283,444)(341,444)(341,281){3}
//: {4}(279,444)(65,444){5}
//: enddecls

  //: joint g4 (w9) @(281, 444) /w:[ 2 1 4 -1 ]
  //: IN g8 (A2) @(3,386) /sn:0 /w:[ 0 ]
  //: joint g13 (A2) @(34, 386) /w:[ 2 -1 1 4 ]
  //: joint g3 (A1) @(149, 355) /w:[ 2 1 4 -1 ]
  _GGAND2 #(6) a3a2_ (.I0(A3), .I1(w7), .Z(w8));   //: @(219,275) /R:1 /w:[ 0 3 0 ]
  //: joint g2 (A3) @(32, 415) /w:[ 1 -1 2 4 ]
  _GGAND2 #(6) a3_a1 (.I0(w9), .I1(A1), .Z(w11));   //: @(284,273) /R:1 /w:[ 0 3 1 ]
  //: joint g1 (w7) @(81, 399) /w:[ 2 4 1 -1 ]
  _GGAND3 #(8) a3_a2a0 (.I0(w9), .I1(A2), .I2(A0), .Z(w14));   //: @(346,270) /R:1 /w:[ 3 3 0 1 ]
  _GGNBUF #(2) g11 (.I(A2), .Z(w7));   //: @(55,399) /sn:0 /w:[ 5 0 ]
  _GGNBUF #(2) g10 (.I(A0), .Z(w1));   //: @(55,337) /sn:0 /w:[ 5 0 ]
  //: IN g6 (A0) @(3,319) /sn:0 /w:[ 3 ]
  //: IN g9 (A3) @(3,415) /sn:0 /w:[ 3 ]
  //: IN g7 (A1) @(3,355) /sn:0 /w:[ 5 ]
  //: OUT g15 (A) @(214,91) /sn:0 /R:1 /w:[ 0 ]
  _GGAND2 #(6) a2_a0_ (.I0(w7), .I1(w1), .Z(w2));   //: @(84,276) /R:1 /w:[ 5 5 1 ]
  //: joint g14 (A0) @(34, 319) /w:[ 1 -1 2 4 ]
  _GGAND2 #(6) a1a0_ (.I0(A1), .I1(w1), .Z(w5));   //: @(152,275) /R:1 /w:[ 0 3 1 ]
  _GGOR5 #(12) g5 (.I0(w2), .I1(w5), .I2(w8), .I3(w11), .I4(w14), .Z(A));   //: @(219,181) /sn:0 /R:1 /w:[ 0 0 1 0 0 1 ]
  //: joint g0 (w1) @(86, 337) /w:[ 2 4 1 -1 ]
  _GGNBUF #(2) g12 (.I(A3), .Z(w9));   //: @(55,444) /sn:0 /w:[ 5 5 ]

endmodule
//: /netlistEnd

//: /netlistBegin segmentoC
module segmentoC(a3, a1, a2, a0, C);
//: interface  /sz:(102, 96) /bd:[ Ri0>a0(16/96) Ri1>a1(32/96) Ri2>a2(48/96) Ri3>a3(64/96) Lo0<C(16/96) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input a2;    //: /sn:0 {0}(473,227)(473,308)(133,308){1}
input a3;    //: /sn:0 {0}(180,328)(133,328){1}
input a1;    //: /sn:0 {0}(180,288)(133,288){1}
input a0;    //: /sn:0 {0}(366,227)(366,268)(133,268){1}
output C;    //: /sn:0 {0}(364,106)(364,61){1}
wire w7;    //: /sn:0 {0}(196,328)(359,328){1}
//: {2}(363,328)(468,328)(468,227){3}
//: {4}(361,326)(361,227){5}
wire w4;    //: /sn:0 {0}(196,288)(261,288)(261,249){1}
//: {2}(261,245)(261,227){3}
//: {4}(259,247)(256,247)(256,227){5}
wire w0;    //: /sn:0 {0}(259,206)(259,142)(359,142)(359,127){1}
wire w3;    //: /sn:0 {0}(471,206)(471,142)(369,142)(369,127){1}
wire w1;    //: /sn:0 {0}(364,206)(364,127){1}
//: enddecls

  //: IN g8 (a3) @(131,328) /sn:0 /w:[ 1 ]
  //: joint g3 (w7) @(361, 328) /w:[ 2 4 1 -1 ]
  //: joint g2 (w4) @(261, 247) /w:[ -1 2 4 1 ]
  _GGNAND3 #(6) g1 (.I0(w0), .I1(w1), .I2(w3), .Z(C));   //: @(364,116) /sn:0 /R:1 /w:[ 1 1 1 0 ]
  _GGNBUF #(2) g11 (.I(a3), .Z(w7));   //: @(186,328) /sn:0 /w:[ 0 0 ]
  _GGNAND2 #(4) a3_a0_ (.I0(w7), .I1(a0), .Z(w1));   //: @(364,216) /R:1 /w:[ 5 0 0 ]
  _GGNBUF #(2) g10 (.I(a1), .Z(w4));   //: @(186,288) /sn:0 /w:[ 0 0 ]
  //: IN g6 (a1) @(131,288) /sn:0 /w:[ 1 ]
  //: IN g7 (a2) @(131,308) /sn:0 /w:[ 1 ]
  _GGNAND2 #(4) a1_ (.I0(w4), .I1(w4), .Z(w0));   //: @(259,216) /R:1 /w:[ 5 3 0 ]
  //: IN g5 (a0) @(131,268) /sn:0 /w:[ 1 ]
  //: OUT g0 (C) @(364,64) /sn:0 /R:1 /w:[ 1 ]
  _GGNAND2 #(4) a3_a2 (.I0(w7), .I1(a2), .Z(w3));   //: @(471,216) /R:1 /w:[ 3 0 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin segmentoG
module segmentoG(a0, a3, a2, G, a1);
//: interface  /sz:(102, 96) /bd:[ Ri0>a0(16/96) Ri1>a1(32/96) Ri2>a2(48/96) Ri3>a3(64/96) Lo0<G(16/96) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input a2;    //: /sn:0 {0}(170,222)(252,222)(252,223)(264,223){1}
input a3;    //: /sn:0 {0}(170,200)(216,200)(216,213)(264,213){1}
output G;    //: /sn:0 {0}(518,160)(487,160){1}
input a1;    //: /sn:0 {0}(170,246)(224,246)(224,233)(264,233){1}
input a0;    //: /sn:0 {0}(366,38)(366,80){1}
supply1 w13;    //: /sn:0 {0}(225,104)(225,153)(264,153){1}
//: {2}(268,153)(299,153){3}
//: {4}(266,151)(266,119)(312,119)(312,129){5}
wire w6;    //: /sn:0 {0}(384,149)(328,149){1}
wire w7;    //: /sn:0 {0}(328,156)(361,156)(361,165)(466,165){1}
wire w4;    //: /sn:0 {0}(328,142)(440,142)(440,155)(466,155){1}
wire w3;    //: /sn:0 {0}(328,136)(451,136)(451,150)(466,150){1}
wire [2:0] w1;    //: /sn:0 {0}(#:270,223)(312,223)(312,175){1}
wire w8;    //: /sn:0 {0}(328,163)(343,163){1}
wire w18;    //: /sn:0 {0}(328,129)(340,129){1}
wire w12;    //: /sn:0 {0}(405,152)(429,152)(429,160)(466,160){1}
wire w2;    //: /sn:0 {0}(384,154)(366,154)(366,96){1}
wire w10;    //: /sn:0 {0}(328,176)(451,176)(451,170)(466,170){1}
wire w9;    //: /sn:0 {0}(328,169)(343,169){1}
//: enddecls

  _GGDEMUX8 #(1, 1, 1) g4 (.F(w13), .S(w1), .E(w13), .Z0(w18), .Z1(w3), .Z2(w4), .Z3(w6), .Z4(w7), .Z5(w8), .Z6(w9), .Z7(w10));   //: @(312,153) /sn:0 /R:1 /w:[ 3 1 5 0 0 0 1 0 0 0 0 ] /ss:0 /do:1
  _GGOR5 #(12) g8 (.I0(w3), .I1(w4), .I2(w12), .I3(w7), .I4(w10), .Z(G));   //: @(477,160) /sn:0 /w:[ 1 1 1 1 1 1 ]
  //: IN g3 (a0) @(366,36) /sn:0 /R:3 /w:[ 0 ]
  //: IN g2 (a3) @(168,200) /sn:0 /w:[ 0 ]
  //: IN g1 (a2) @(168,222) /sn:0 /w:[ 0 ]
  //: OUT g11 (G) @(515,160) /sn:0 /w:[ 0 ]
  _GGAND2 #(6) g10 (.I0(w6), .I1(w2), .Z(w12));   //: @(395,152) /sn:0 /w:[ 0 0 0 ]
  //: VDD g6 (w13) @(236,104) /sn:0 /w:[ 0 ]
  //: joint g7 (w13) @(266, 153) /w:[ 2 4 1 -1 ]
  _GGNBUF #(2) g9 (.I(a0), .Z(w2));   //: @(366,86) /sn:0 /R:3 /w:[ 1 1 ]
  assign w1 = {a3, a2, a1}; //: CONCAT g5  @(269,223) /sn:0 /w:[ 0 1 1 1 ] /dr:0 /tp:0 /drp:1
  //: IN g0 (a1) @(168,246) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin segmentoB
module segmentoB(B, a3, a2, a1, a0);
//: interface  /sz:(160, 96) /bd:[ Ti0>a0(20/160) Ti1>a1(60/160) Ti2>a2(100/160) Ti3>a3(140/160) Lo0<B(46/96) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output B;    //: /sn:0 {0}(452,66)(452,29){1}
input a2;    //: /sn:0 {0}(192,352)(234,352){1}
input a3;    //: /sn:0 {0}(191,389)(233,389){1}
input a1;    //: /sn:0 {0}(356,190)(356,276)(212,276){1}
//: {2}(208,276)(192,276){3}
//: {4}(210,278)(210,315)(234,315){5}
input a0;    //: /sn:0 {0}(234,255)(212,255)(212,228){1}
//: {2}(214,226)(457,226)(457,190){3}
//: {4}(210,226)(192,226){5}
wire w7;    //: /sn:0 {0}(540,190)(540,389)(249,389){1}
wire w4;    //: /sn:0 {0}(452,190)(452,313){1}
//: {2}(454,315)(545,315)(545,190){3}
//: {4}(450,315)(250,315){5}
wire w0;    //: /sn:0 {0}(351,190)(351,350){1}
//: {2}(353,352)(447,352)(447,190){3}
//: {4}(349,352)(250,352){5}
wire w1;    //: /sn:0 {0}(250,255)(361,255)(361,190){1}
wire w2;    //: /sn:0 {0}(447,87)(447,102)(356,102)(356,169){1}
wire w10;    //: /sn:0 {0}(542,169)(542,102)(457,102)(457,87){1}
wire w5;    //: /sn:0 {0}(452,87)(452,169){1}
//: enddecls

  //: joint g8 (w0) @(351, 352) /w:[ 2 1 4 -1 ]
  _GGNBUF #(2) g4 (.I(a0), .Z(w1));   //: @(240,255) /sn:0 /w:[ 0 0 ]
  //: OUT g13 (B) @(452,32) /sn:0 /R:1 /w:[ 1 ]
  //: IN g3 (a3) @(189,389) /sn:0 /w:[ 0 ]
  //: IN g2 (a2) @(190,352) /sn:0 /w:[ 0 ]
  //: IN g1 (a1) @(190,276) /sn:0 /w:[ 3 ]
  //: joint g11 (w4) @(452, 315) /w:[ 2 1 4 -1 ]
  _GGOR3 #(8) a2_a1_a0 (.I0(w0), .I1(w4), .I2(a0), .Z(w5));   //: @(452,179) /R:1 /w:[ 3 0 3 1 ]
  _GGOR2 #(6) a3_a1_ (.I0(w7), .I1(w4), .Z(w10));   //: @(542,179) /R:1 /w:[ 0 3 0 ]
  //: joint g10 (a0) @(212, 226) /w:[ 2 -1 4 1 ]
  _GGNBUF #(2) g6 (.I(a2), .Z(w0));   //: @(240,352) /sn:0 /w:[ 1 5 ]
  //: joint g9 (a1) @(210, 276) /w:[ 1 -1 2 4 ]
  _GGNBUF #(2) g7 (.I(a3), .Z(w7));   //: @(239,389) /sn:0 /w:[ 1 1 ]
  _GGNBUF #(2) g5 (.I(a1), .Z(w4));   //: @(240,315) /sn:0 /w:[ 5 5 ]
  _GGOR3 #(8) a2_a1a0_ (.I0(w0), .I1(a1), .I2(w1), .Z(w2));   //: @(356,179) /R:1 /w:[ 0 0 1 1 ]
  //: IN g0 (a0) @(190,226) /sn:0 /w:[ 5 ]
  _GGAND3 #(8) g12 (.I0(w2), .I1(w5), .I2(w10), .Z(B));   //: @(452,76) /sn:0 /R:1 /w:[ 0 0 1 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin segmentoD
module segmentoD(a2, a1, a0, a3, D);
//: interface  /sz:(102, 80) /bd:[ Ri0>a0(16/80) Ri1>a1(32/80) Ri2>a2(48/80) Ri3>a3(64/80) To0<D(20/102) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input a2;    //: /sn:0 {0}(113,390)(80,390)(80,354){1}
//: {2}(82,352)(626,352)(626,187){3}
//: {4}(78,352)(65,352){5}
input a3;    //: /sn:0 {0}(621,187)(621,423)(65,423){1}
input a1;    //: /sn:0 {0}(631,187)(631,289)(386,289){1}
//: {2}(384,287)(384,187){3}
//: {4}(382,289)(88,289){5}
//: {6}(84,289)(65,289){7}
//: {8}(86,291)(86,318)(113,318){9}
input a0;    //: /sn:0 {0}(65,234)(84,234){1}
//: {2}(88,234)(389,234)(389,187){3}
//: {4}(86,236)(86,260)(113,260){5}
output D;    //: /sn:0 {0}(516,47)(516,95){1}
wire w0;    //: /sn:0 {0}(511,116)(511,131)(384,131)(384,166){1}
wire w3;    //: /sn:0 {0}(628,166)(628,131)(521,131)(521,116){1}
wire w1;    //: /sn:0 {0}(516,167)(516,116){1}
wire w8;    //: /sn:0 {0}(516,188)(516,318)(129,318){1}
wire w2;    //: /sn:0 {0}(379,187)(379,388){1}
//: {2}(381,390)(511,390)(511,188){3}
//: {4}(377,390)(129,390){5}
wire w9;    //: /sn:0 {0}(636,187)(636,260)(523,260){1}
//: {2}(521,258)(521,188){3}
//: {4}(519,260)(129,260){5}
//: enddecls

  //: IN g4 (a2) @(63,352) /sn:0 /w:[ 5 ]
  _GGNBUF #(2) g8 (.I(a2), .Z(w2));   //: @(119,390) /sn:0 /w:[ 0 5 ]
  //: IN g3 (a1) @(63,289) /sn:0 /w:[ 7 ]
  //: joint g13 (a1) @(384, 289) /w:[ 1 2 4 -1 ]
  //: IN g2 (a0) @(63,234) /sn:0 /w:[ 0 ]
  _GGNOR3 #(6) g1 (.I0(w0), .I1(w1), .I2(w3), .Z(D));   //: @(516,105) /sn:0 /R:1 /w:[ 0 1 1 1 ]
  //: joint g11 (a0) @(86, 234) /w:[ 2 -1 1 4 ]
  //: joint g10 (a1) @(86, 289) /w:[ 5 -1 6 8 ]
  _GGNBUF #(2) g6 (.I(a0), .Z(w9));   //: @(119,260) /sn:0 /w:[ 5 5 ]
  _GGNBUF #(2) g7 (.I(a1), .Z(w8));   //: @(119,318) /sn:0 /w:[ 9 1 ]
  //: joint g9 (w2) @(379, 390) /w:[ 2 1 4 -1 ]
  _GGNOR4 #(8) a3a2a1a0_ (.I0(a3), .I1(a2), .I2(a1), .I3(w9), .Z(w3));   //: @(628,176) /R:1 /w:[ 0 3 0 0 0 ]
  //: IN g5 (a3) @(63,423) /sn:0 /w:[ 1 ]
  //: joint g14 (w9) @(521, 260) /w:[ 1 2 4 -1 ]
  //: OUT g0 (D) @(516,50) /sn:0 /R:1 /w:[ 0 ]
  _GGNOR3 #(6) a2_a1_a0_ (.I0(w2), .I1(w8), .I2(w9), .Z(w1));   //: @(516,177) /R:1 /w:[ 3 0 3 0 ]
  //: joint g12 (a2) @(80, 352) /w:[ 2 -1 4 1 ]
  _GGNOR3 #(6) a2_a1a0 (.I0(w2), .I1(a1), .I2(a0), .Z(w0));   //: @(384,176) /R:1 /w:[ 0 3 3 1 ]

endmodule
//: /netlistEnd

//: /netlistBegin segmentoE
module segmentoE(E, a2, a1, a0, a3);
//: interface  /sz:(160, 80) /bd:[ Bi0>a0(20/160) Bi1>a1(60/160) Bi2>a2(100/160) Bi3>a3(140/160) Ro0<E(16/80) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
supply1 w6;    //: /sn:0 {0}(250,170)(145,170)(145,159){1}
//: {2}(147,157)(250,157){3}
//: {4}(145,155)(145,146){5}
//: {6}(147,144)(250,144){7}
//: {8}(145,142)(145,49){9}
input a2;    //: /sn:0 {0}(204,59)(204,92){1}
input a3;    //: /sn:0 {0}(249,271)(249,240)(256,240)(256,225){1}
input a1;    //: /sn:0 {0}(266,269)(266,225){1}
input a0;    //: /sn:0 {0}(290,271)(290,240)(276,240)(276,225){1}
output E;    //: /sn:0 {0}(279,154)(306,154)(306,155)(334,155){1}
supply0 w5;    //: /sn:0 {0}(250,177)(179,177){1}
//: {2}(177,175)(177,166){3}
//: {4}(179,164)(250,164){5}
//: {6}(177,162)(177,152){7}
//: {8}(179,150)(250,150){9}
//: {10}(177,148)(177,137)(250,137){11}
//: {12}(177,179)(177,218){13}
wire [2:0] w15;    //: /sn:0 {0}(#:266,219)(266,177){1}
wire w1;    //: /sn:0 {0}(204,108)(204,130)(250,130){1}
//: enddecls

  _GGMUX8 #(20, 20) g4 (.I0(w1), .I1(w5), .I2(w6), .I3(w5), .I4(w6), .I5(w5), .I6(w6), .I7(w5), .S(w15), .Z(E));   //: @(266,154) /sn:0 /R:1 /w:[ 1 11 7 9 3 5 0 0 1 0 ] /ss:0 /do:1
  //: joint g8 (w5) @(177, 177) /w:[ 1 2 -1 12 ]
  //: VDD g3 (w6) @(156,49) /sn:0 /w:[ 9 ]
  //: joint g13 (w6) @(145, 144) /w:[ 6 8 -1 5 ]
  //: GROUND g2 (w5) @(177,224) /sn:0 /w:[ 13 ]
  //: OUT g1 (E) @(331,155) /sn:0 /w:[ 1 ]
  //: IN g11 (a2) @(204,57) /sn:0 /R:3 /w:[ 0 ]
  //: joint g10 (w5) @(177, 164) /w:[ 4 6 -1 3 ]
  //: IN g6 (a1) @(266,271) /sn:0 /R:1 /w:[ 0 ]
  //: IN g7 (a0) @(290,273) /sn:0 /R:1 /w:[ 0 ]
  //: joint g9 (w6) @(145, 157) /w:[ 2 4 -1 1 ]
  //: IN g5 (a3) @(249,273) /sn:0 /R:1 /w:[ 0 ]
  //: joint g14 (w5) @(177, 150) /w:[ 8 10 -1 7 ]
  assign w15 = {a3, a1, a0}; //: CONCAT g0  @(266,220) /sn:0 /R:1 /w:[ 0 1 1 1 ] /dr:0 /tp:1 /drp:1
  _GGNBUF #(2) g12 (.I(a2), .Z(w1));   //: @(204,98) /sn:0 /R:3 /w:[ 1 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin segmentoF
module segmentoF(a2, a0, a1, E, a3);
//: interface  /sz:(160, 80) /bd:[ Bi0>a3(140/160) Bi1>a2(100/160) Bi2>a1(60/160) Bi3>a0(20/160) Ro0<E(59/80) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input a2;    //: /sn:0 {0}(153,229)(114,229)(114,239)(58,239){1}
input a3;    //: /sn:0 {0}(57,219)(153,219){1}
input a1;    //: /sn:0 {0}(58,269)(137,269)(137,239)(153,239){1}
input a0;    //: /sn:0 {0}(305,44)(305,-5){1}
supply1 w10;    //: /sn:0 {0}(219,161)(219,205){1}
output E;    //: /sn:0 {0}(481,220)(523,220)(523,209)(612,209){1}
wire w6;    //: /sn:0 {0}(235,232)(370,232)(370,223)(460,223){1}
wire w7;    //: /sn:0 {0}(235,238)(250,238){1}
wire w16;    //: /sn:0 {0}(396,262)(445,262)(445,233)(460,233){1}
wire w4;    //: /sn:0 {0}(235,218)(445,218)(445,213)(460,213){1}
wire w15;    //: /sn:0 {0}(235,245)(381,245)(381,228)(460,228){1}
wire [2:0] w0;    //: /sn:0 {0}(#:159,229)(206,229){1}
wire w3;    //: /sn:0 {0}(235,212)(250,212){1}
wire w1;    //: /sn:0 {0}(399,127)(450,127)(450,208)(460,208){1}
wire w17;    //: /sn:0 {0}(378,129)(290,129)(290,205)(235,205){1}
wire w11;    //: /sn:0 {0}(378,124)(363,124)(363,122)(307,122){1}
//: {2}(305,120)(305,60){3}
//: {4}(305,124)(305,154){5}
//: {6}(307,156)(377,156){7}
//: {8}(305,158)(305,259)(375,259){9}
wire w13;    //: /sn:0 {0}(398,159)(445,159)(445,218)(460,218){1}
wire w5;    //: /sn:0 {0}(235,225)(363,225)(363,161)(377,161){1}
wire w9;    //: /sn:0 {0}(375,264)(251,264)(251,252)(235,252){1}
//: enddecls

  //: IN g4 (a2) @(56,239) /sn:0 /w:[ 1 ]
  //: IN g8 (a0) @(305,-7) /sn:0 /R:3 /w:[ 1 ]
  _GGAND2 #(6) g13 (.I0(w11), .I1(w9), .Z(w16));   //: @(386,262) /sn:0 /w:[ 9 0 0 ]
  //: IN g3 (a1) @(56,269) /sn:0 /w:[ 0 ]
  assign w0 = {a3, a2, a1}; //: CONCAT g2  @(158,229) /sn:0 /w:[ 0 1 0 1 ] /dr:0 /tp:1 /drp:1
  //: VDD g1 (w10) @(230,161) /sn:0 /w:[ 0 ]
  _GGAND2 #(6) g11 (.I0(w11), .I1(w17), .Z(w1));   //: @(389,127) /sn:0 /w:[ 0 0 0 ]
  _GGNBUF #(2) g10 (.I(a0), .Z(w11));   //: @(305,50) /sn:0 /R:3 /w:[ 0 3 ]
  //: OUT g6 (E) @(609,209) /sn:0 /w:[ 1 ]
  _GGAND2 #(6) g9 (.I0(w11), .I1(w5), .Z(w13));   //: @(388,159) /sn:0 /w:[ 7 1 0 ]
  _GGOR6 #(14) g7 (.I0(w1), .I1(w4), .I2(w13), .I3(w6), .I4(w15), .I5(w16), .Z(E));   //: @(471,220) /sn:0 /w:[ 1 1 1 1 1 1 0 ]
  //: joint g14 (w11) @(305, 156) /w:[ 6 5 -1 8 ]
  //: IN g5 (a3) @(55,219) /sn:0 /w:[ 0 ]
  _GGDECODER8 #(6, 6) g0 (.I(w0), .E(w10), .Z0(w17), .Z1(w3), .Z2(w4), .Z3(w5), .Z4(w6), .Z5(w7), .Z6(w15), .Z7(w9));   //: @(219,229) /sn:0 /R:1 /w:[ 1 1 1 0 0 0 0 0 0 1 ] /ss:1 /do:1
  //: joint g12 (w11) @(305, 122) /w:[ 1 2 -1 4 ]

endmodule
//: /netlistEnd

